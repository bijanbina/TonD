test1

V1 1 0 1
V2 2 7 DC 0 $ <---- ammeter
R1 7 1 5
R2 3 0 10
E1 2 0 3 0 2
V3 3 4 DC 0 $ <---- output
L1 4 1 0.5 IC=0
F1 3 2 v2 2
 

.control
	TRAN	0.1us 2ms
.endc

.end
